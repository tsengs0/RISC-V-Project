module RegFile (
	input wire []
);
