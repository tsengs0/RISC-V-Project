`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Bo-Yu Tseng
// 
// Create Date: 04.Jan.2023
// Design: rv32_core
// Project Name: RISC-V core IP development
// Target Devices: Xilinx FPGAs and open source ASIC process
// Tool Versions: 
// Description: 
// 				A RTL module of instruction decoder for RV32I
// Dependencies: 
// 				a) ../macros/rv32_define.vh
//				b) ../macros/define.vh
// Revision:
// Additional Comments:
//     
//////////////////////////////////////////////////////////////////////////////////
